// platform.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module platform (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

endmodule
